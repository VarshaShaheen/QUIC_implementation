`timescale 1ns/10ps

module tb;

reg clk;
reg encoded;
wire [463:0] decoded;
wire [15:0] source_port;
wire [15:0] dest_port;
wire [133:0] data;

integer i;

// Instantiate the design under test
pass_through dut (
    .clk(clk),
    .encoded(encoded),
    .decoded(decoded),
    .source_port(source_port),
    .dest_port(dest_port),
    .data(data)
);

// Clock generation
always begin
    #5 clk = ~clk;
end

// Define Ethernet frame
localparam ETH_FRAME_LEN = 976;
reg [ETH_FRAME_LEN-1:0] eth_frame = 976'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010011010101010101010101010100110101001100110101010101010101010101010101010101001100110010110101010101010101010101010101010100110101010101010101010101010101001101010101010101010011010100101100101100101011001011001011010010110101010101001100110011010101010101010101001101010101010011001011010101010100110011001101010101010101010100110101010101001011010100101010101100110101010101010101001010101011001101010101001101010101010101010101001100101011010101010101010101010101010101010011010011010101001011010011001100101100101101010010110010110101001011001010101101001101010101010011001100101011001011001010101100101011010011010010110010110101001011010011010
10100110101010101010011010101001101001101010100110100110101010010101010101010101101010101001101010101010010101101010010110101010;

initial begin
    // Initialize inputs
    clk = 0;
    encoded = 0;

    // Apply Ethernet frame to encoded input bit by bit
    for (i = 0; i < ETH_FRAME_LEN; i = i+1) begin
        @(posedge clk);
        encoded = eth_frame[i];
    end
    
    encoded = 0;

    // Check outputs
    // ...
end

endmodule
